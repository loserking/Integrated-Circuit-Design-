`timescale 1ns/1ps

module DOQE_ppl(clk,rst,A,B,C,D,DOQE_ppl_num);
// DO NOT CHANGE !
	input			clk;
	input			rst;
	input		[3:0]	A;
	input		[6:0]	B;
	input   [5:0] C;
	
	output	[14:0]D;
    output  [50:0]  DOQE_ppl_num;	

  // Write your design here


endmodule

