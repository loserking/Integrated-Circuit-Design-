`timescale 1ns/1ps
module COMPARATOR_51(min, i0, i1, i2, i3, i4);
	//DO NOT CHANGE!
	output [2:0] min;
	input  [5:0] i0, i1, i2, i3, i4;
	
	//---------------------------------------------------
	//Write your design here




endmodule 